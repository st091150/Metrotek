
module const_ffff(
    output [15:0] result
);
    assign result = 16'hFFFF;
endmodule


module const_A001(
    output [15:0] result
);
    assign result = 16'hA001;
endmodule
