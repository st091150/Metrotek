
module const_ffff(
    output [15:0] result
);
    assign result = 16'hFFFF;
endmodule


module const_8005(
    output [15:0] result
);
    assign result = 16'h8005;
endmodule
