// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details.

// PROGRAM		"Quartus Prime"
// VERSION		"Version 18.1.0 Build 625 09/12/2018 SJ Lite Edition"
// CREATED		"Tue Nov  4 02:57:26 2025"

module mux161 (
	GN,
	IN12,
	IN13,
	IN14,
	IN15,
	IN4,
	IN5,
	IN6,
	IN7,
	IN8,
	IN9,
	IN10,
	IN11,
	SEL2,
	SEL1,
	SEL0,
	SEL3,
	IN0,
	IN1,
	IN2,
	IN3,
	OUT1
);


input wire	GN;
input wire	IN12;
input wire	IN13;
input wire	IN14;
input wire	IN15;
input wire	IN4;
input wire	IN5;
input wire	IN6;
input wire	IN7;
input wire	IN8;
input wire	IN9;
input wire	IN10;
input wire	IN11;
input wire	SEL2;
input wire	SEL1;
input wire	SEL0;
input wire	SEL3;
input wire	IN0;
input wire	IN1;
input wire	IN2;
input wire	IN3;
output wire	OUT1;

wire	SYNTHESIZED_WIRE_88;
wire	SYNTHESIZED_WIRE_89;
wire	SYNTHESIZED_WIRE_90;
wire	SYNTHESIZED_WIRE_91;
wire	SYNTHESIZED_WIRE_92;
wire	SYNTHESIZED_WIRE_93;
wire	SYNTHESIZED_WIRE_94;
wire	SYNTHESIZED_WIRE_34;
wire	SYNTHESIZED_WIRE_35;
wire	SYNTHESIZED_WIRE_36;
wire	SYNTHESIZED_WIRE_37;
wire	SYNTHESIZED_WIRE_38;
wire	SYNTHESIZED_WIRE_39;
wire	SYNTHESIZED_WIRE_40;
wire	SYNTHESIZED_WIRE_41;
wire	SYNTHESIZED_WIRE_42;
wire	SYNTHESIZED_WIRE_43;
wire	SYNTHESIZED_WIRE_44;
wire	SYNTHESIZED_WIRE_45;
wire	SYNTHESIZED_WIRE_46;
wire	SYNTHESIZED_WIRE_47;
wire	SYNTHESIZED_WIRE_48;
wire	SYNTHESIZED_WIRE_49;
wire	SYNTHESIZED_WIRE_95;
wire	SYNTHESIZED_WIRE_53;
wire	SYNTHESIZED_WIRE_96;
wire	SYNTHESIZED_WIRE_57;
wire	SYNTHESIZED_WIRE_58;
wire	SYNTHESIZED_WIRE_59;
wire	SYNTHESIZED_WIRE_60;
wire	SYNTHESIZED_WIRE_61;
wire	SYNTHESIZED_WIRE_74;
wire	SYNTHESIZED_WIRE_78;




assign	SYNTHESIZED_WIRE_41 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_90 & IN9;

assign	SYNTHESIZED_WIRE_93 =  ~SEL0;

assign	SYNTHESIZED_WIRE_91 =  ~SEL2;

assign	SYNTHESIZED_WIRE_95 =  ~SYNTHESIZED_WIRE_91;

assign	SYNTHESIZED_WIRE_92 =  ~SEL3;

assign	SYNTHESIZED_WIRE_96 =  ~SYNTHESIZED_WIRE_92;

assign	SYNTHESIZED_WIRE_88 =  ~GN;

assign	SYNTHESIZED_WIRE_90 =  ~SYNTHESIZED_WIRE_93;

assign	SYNTHESIZED_WIRE_89 =  ~SEL1;

assign	SYNTHESIZED_WIRE_94 =  ~SYNTHESIZED_WIRE_89;

assign	SYNTHESIZED_WIRE_49 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_90 & IN1;

assign	SYNTHESIZED_WIRE_48 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_94 & SYNTHESIZED_WIRE_90 & IN3;

assign	SYNTHESIZED_WIRE_45 = IN5 & SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_90 & SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_44 = IN7 & SYNTHESIZED_WIRE_94 & SYNTHESIZED_WIRE_90 & SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_38 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_93 & IN8;

assign	SYNTHESIZED_WIRE_40 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_94 & SYNTHESIZED_WIRE_90 & IN11;

assign	SYNTHESIZED_WIRE_34 = IN12 & SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_93 & SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_37 = IN13 & SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_90 & SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_36 = IN15 & SYNTHESIZED_WIRE_94 & SYNTHESIZED_WIRE_90 & SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_57 = SYNTHESIZED_WIRE_34 | SYNTHESIZED_WIRE_35 | SYNTHESIZED_WIRE_36 | SYNTHESIZED_WIRE_37;

assign	SYNTHESIZED_WIRE_78 = SYNTHESIZED_WIRE_38 | SYNTHESIZED_WIRE_39 | SYNTHESIZED_WIRE_40 | SYNTHESIZED_WIRE_41;

assign	SYNTHESIZED_WIRE_53 = SYNTHESIZED_WIRE_42 | SYNTHESIZED_WIRE_43 | SYNTHESIZED_WIRE_44 | SYNTHESIZED_WIRE_45;

assign	SYNTHESIZED_WIRE_74 = SYNTHESIZED_WIRE_46 | SYNTHESIZED_WIRE_47 | SYNTHESIZED_WIRE_48 | SYNTHESIZED_WIRE_49;

assign	SYNTHESIZED_WIRE_61 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_92 & SYNTHESIZED_WIRE_95 & SYNTHESIZED_WIRE_53;

assign	SYNTHESIZED_WIRE_60 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_96 & SYNTHESIZED_WIRE_95 & SYNTHESIZED_WIRE_57;

assign	OUT1 = SYNTHESIZED_WIRE_58 | SYNTHESIZED_WIRE_59 | SYNTHESIZED_WIRE_60 | SYNTHESIZED_WIRE_61;

assign	SYNTHESIZED_WIRE_46 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_93 & IN0;

assign	SYNTHESIZED_WIRE_39 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_94 & SYNTHESIZED_WIRE_93 & IN10;

assign	SYNTHESIZED_WIRE_35 = IN14 & SYNTHESIZED_WIRE_94 & SYNTHESIZED_WIRE_93 & SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_58 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_92 & SYNTHESIZED_WIRE_91 & SYNTHESIZED_WIRE_74;

assign	SYNTHESIZED_WIRE_59 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_96 & SYNTHESIZED_WIRE_91 & SYNTHESIZED_WIRE_78;

assign	SYNTHESIZED_WIRE_47 = SYNTHESIZED_WIRE_88 & SYNTHESIZED_WIRE_94 & SYNTHESIZED_WIRE_93 & IN2;

assign	SYNTHESIZED_WIRE_42 = IN4 & SYNTHESIZED_WIRE_89 & SYNTHESIZED_WIRE_93 & SYNTHESIZED_WIRE_88;

assign	SYNTHESIZED_WIRE_43 = IN6 & SYNTHESIZED_WIRE_94 & SYNTHESIZED_WIRE_93 & SYNTHESIZED_WIRE_88;


endmodule
